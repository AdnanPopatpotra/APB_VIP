/* -.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.

* Company       : SCALEDGE
* Created By    : MOHAMADADNAN POPATPOTRA
* File Name 	: apb_simple_read_tc.sv
* Creation Date : 02-08-2023
* Last Modified : 02-08-2023 12:05:57
* Purpose       :  
_._._._._._._._._._._._._._._._._._._._._.*/


