/* -.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.

* Company       : SCALEDGE
* Created By    : MOHAMADADNAN POPATPOTRA
* File Name 	: apb_defines.sv
* Creation Date : 24-07-2023
* Last Modified : 31-08-2023 15:10:51
* Purpose       :  
_._._._._._._._._._._._._._._._._._._._._.*/

`ifndef APB_DEFINES_SV
`define APB_DEFINES_SV

`define ADDR_WIDTH 5
`define DATA_WIDTH 8
`define TIMEOUT 20

`endif
